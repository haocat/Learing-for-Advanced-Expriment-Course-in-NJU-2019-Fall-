`timescale 1ns / 1ps
module simu2(

    );
     parameter k=484;
       parameter n=511;
       reg clk;
       reg rst;
       reg [k-1:0]msg;
       reg [3:0]send;
       wire [n-1:0]bch_dataout;
       reg [8:0]i=484;
       always #5 clk = ~clk;
       
       initial
       begin
           msg[k-1:0]=484'b1101100111011010011110111110101000011010001100011101100010101011111000101010001001111011010011101000010101011100010111000101110001010000111011010000000011000100100000111000100011101010100110110000111110110111110000100000010011000010110000010010110100111001100101110001010101111010011011111100100011100100101110111110010000110010110001000000110100110101111100100111000101100000100100101110101110100000001011100011011110011000000101111101011000110110101000010100010001010101000111011111;
           clk=1;
           rst=1;
           #102 rst=~rst;
         /*               send[3]<=msg[i-1];
             send[2]<=msg[i-2];
             send[1]<=msg[i-3];
             send[0]<=msg[i-4];
             i = i-4;*/
       end    
       
        always @(negedge clk)
        begin
           if (i>3&&!rst&&i)
               begin 
               send[3]<=msg[i-1];
               send[2]<=msg[i-2];
               send[1]<=msg[i-3];
               send[0]<=msg[i-4];
               i = i-4;
               end
       end
               
       pa1 out(
           .rst(rst),
           .clk(clk),
           .msg(send),
           .bch_dataout(bch_dataout)
           );
endmodule
